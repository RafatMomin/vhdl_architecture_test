library IEEE;
use IEEE.std_logic_1164.all;

entity reg_nbit is
  generic (N : integer := 32); -- Number of bits
  port (
    i_CLK  : in std_logic;     -- Clock input
    i_RST  : in std_logic;     -- Reset input
    i_WE   : in std_logic;     -- Write enable input
    i_D    : in std_logic_vector(N-1 downto 0); -- Data input
    o_Q    : out std_logic_vector(N-1 downto 0) -- Data output
  );
end reg_nbit;

architecture structural of reg_nbit is
  component dffg
    port (
      i_CLK  : in std_logic;    
      i_RST  : in std_logic;     
      i_WE   : in std_logic;     
      i_D    : in std_logic;     
      o_Q    : out std_logic    
    );
  end component;

  signal s_Q : std_logic_vector(N-1 downto 0);

begin
  -- Instantiate N D flip-flops
  gen: for i in 0 to N-1 generate
    FF: dffg
      port map(
        i_CLK => i_CLK,
        i_RST => i_RST,
        i_WE  => i_WE,
        i_D   => i_D(i),
        o_Q   => s_Q(i)
      );
  end generate;

  -- Output
  o_Q <= s_Q;

end structural;

